package cover_enable_pkg;

    typedef enum bit {COV_ENABLE, COV_DISABLE} cover_e;
    
endpackage